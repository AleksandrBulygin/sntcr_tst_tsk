
module clockDecrease (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
